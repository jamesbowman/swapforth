`timescale 1 ns / 1 ps

`default_nettype none
`define WIDTH 16

// module progmem #(
//     parameter DATA = 16,
//     parameter ADDR = 3
// ) (
//     input   wire                clk,
//     input   wire    [ADDR-1:0]  addr,
//     // input   wire                wr,
//     // input   wire    [DATA-1:0]  din,
//     output  reg     [DATA-1:0]  dout
// );
//  
//   reg [DATA-1:0] mem [(2**ADDR)-1:0];
//   initial begin
//     $readmemh("compiler/build/nuc.hex", mem);
//   end
//  
//   always @(posedge clk) begin
//     dout      <= mem[addr];
//   end
// endmodule

// module bootrom (
//     input   wire           clk,
//     input   wire    [2:0]  addr,
//     output  reg     [15:0] dout
// );
//   always @(posedge clk)
//     case (addr)
// `include "compiler/build/nuc.v"
//     endcase
// 
// endmodule

module test (
        input clk, we,
        input [7:0] addr,
        input [7:0] wdata,
        output reg [7:0] rdata
);
        reg [7:0] mem [0:255];
        // initial $readmemh("compiler/build/foo.hex", mem);
        always @(posedge clk) begin
                if (we)
                        mem[addr] <= wdata;
                rdata <= mem[addr];
        end
endmodule

module SB_RAM2048x2(
	output [1:0] RDATA,
	input        RCLK, RCLKE, RE,
	input  [10:0] RADDR,
	input         WCLK, WCLKE, WE,
	input  [10:0] WADDR,
	input  [1:0] MASK, WDATA
);
	parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
	parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

  wire [15:0] rd;

  SB_RAM40_4K #(
    .WRITE_MODE(3),
    .READ_MODE(3),
    .INIT_0(INIT_0),
    .INIT_1(INIT_1),
    .INIT_2(INIT_2),
    .INIT_3(INIT_3),
    .INIT_4(INIT_4),
    .INIT_5(INIT_5),
    .INIT_6(INIT_6),
    .INIT_7(INIT_7),
    .INIT_8(INIT_8),
    .INIT_9(INIT_9),
    .INIT_A(INIT_A),
    .INIT_B(INIT_B),
    .INIT_C(INIT_C),
    .INIT_D(INIT_D),
    .INIT_E(INIT_E),
    .INIT_F(INIT_F)
  ) _ram (
    .RDATA(rd),
    .RADDR(RADDR),
    .RCLK(RCLK), .RCLKE(RCLKE), .RE(RE),
    .WCLK(WCLK), .WCLKE(WCLKE), .WE(WE),
    .WADDR(WADDR),
    .MASK(16'h0000), .WDATA({4'b0, WDATA[1], 7'b0, WDATA[0], 3'b0}));

  assign RDATA[0] = rd[3];
  assign RDATA[1] = rd[11];

endmodule

module top(input clk, output D1, output D2, output D3, output D4, output D5,
           output TXD,
           input RXD,
           input resetq,
           output J3_10
);
  localparam MHZ = 12;

  wire io_rd, io_wr;
  wire [15:0] mem_din;
  wire [15:0] mem_addr;
  wire mem_wr;
  wire [15:0] dout;
  wire [15:0] io_din;
  wire [12:0] code_addr;

  wire [15:0] insn;
  reg unlocked = 0;

`include "../build/ram.v"

  j1 _j1(
    .clk(clk),
    .resetq(resetq),
    .io_rd(io_rd),
    .io_wr(io_wr),
    .mem_wr(mem_wr),
    .dout(dout),
    .io_din(io_din),
    .mem_din(mem_din),
    .mem_addr(mem_addr),
    .code_addr(code_addr),
    .insn(insn));

  reg  io_wr_, io_rd_;
  reg [15:0] dout_;
  reg [1:0] io_addr_;

  always @(posedge clk) begin
    {io_rd_, io_wr_, dout_} <= {io_rd, io_wr, dout};
    if (io_rd | io_wr)
      io_addr_ <= mem_addr[1:0];
  end

  assign J3_10 = io_wr;

  wire uart0_valid, uart0_busy;
  wire [7:0] uart0_data;
  wire uart0_wr = io_wr_ & (io_addr_ == 2'b1);
  wire uart0_rd = io_rd_ & (io_addr_ == 2'b1);
  reg [31:0] uart_baud = 32'd115200;
  wire UART0_RX;
  buart #(.CLKFREQ(MHZ * 1000000)) _uart0 (
     .clk(clk),
     .resetq(1'b1),
     .baud(uart_baud),
     .rx(RXD),
     .tx(TXD),
     .rd(uart0_rd),
     .wr(uart0_wr),
     .valid(uart0_valid),
     .busy(uart0_busy),
     .tx_data(dout_[7:0]),
     .rx_data(uart0_data));

  assign io_din = io_addr_[0] ? (uart0_valid ? {8'h01, uart0_data} : {16'h0000}) : {15'd0, !uart0_busy};

  reg [4:0] LEDS;
  assign {D1,D2,D3,D4,D5} = LEDS;
  always @(posedge clk)
    if (io_wr_)
      case (io_addr_)
      2'd2: LEDS <= dout_[4:0];
      endcase

  always @(negedge resetq or posedge clk)
    if (!resetq)
      unlocked <= 0;
    else
      unlocked <= unlocked | io_wr_;

endmodule // top
